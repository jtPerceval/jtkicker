/*  This file is part of JTKICKER.
    JTKICKER program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JTKICKER program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JTKICKER.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 11-11-2021 */

module jtsbaskt_snd(
    input               rst,
    input               clk,
    input               snd_cen,    // 3.5MHz
    input               psg_cen,    // 1.7MHz
    // ROM
    output      [12:0]  rom_addr,
    output reg          rom_cs,
    input       [ 7:0]  rom_data,
    input               rom_ok,
    // From main CPU
    input       [ 7:0]  main_dout,
    input               m2s_data,
    input               m2s_on,
    // Sound
    output     [15:0]   pcm_addr,
    input      [ 7:0]   pcm_data,
    input               pcm_ok,

    output signed [15:0] snd,
    output               sample,
    output               peak
);

localparam CNTW=11;

reg  [ 7:0] latch, psg_data, vlm_data, din, rdac;
wire [ 7:0] ram_dout, vlm_mux, dout;
wire        irq_ack, int_n;
wire [ 2:0] pcm_nc;
wire        vlm_ceng, vlm_me_b;
wire [10:0] psg_snd;
reg         ram_cs;
wire        mreq_n, iorq_n, m1_n;
wire [15:0] A;
reg  [ 2:0] snd_en;
wire        rdy1;
reg         vlm_rst, vlm_st, vlm_sel;
wire        vlm_bsy;
reg         psgdata_cs, vlm_data_cs, vlm_ctrl_cs;
reg         latch_cs, cnt_cs, rdac_cs, psg_cs;
reg [CNTW-1:0] cnt;
wire signed
         [9:0] vlm_snd;

assign vlm_mux = ~vlm_sel ? vlm_data :
               ~vlm_me_b ? pcm_data : 8'hff;
assign pcm_addr[15:13]=0;
assign irq_ack = ~iorq_n & ~m1_n;
assign vlm_ceng = snd_cen & ( vlm_me_b | pcm_ok );
assign rom_addr = A[12:0];
assign sample   = psg_cen;

always @(posedge clk, posedge rst) begin
    if( rst ) begin
        latch    <= 0;
        psg_data <= 0;
        cnt      <= 0;
        snd_en   <= 0;
        vlm_rst  <= 1;
        vlm_st   <= 0;
        vlm_sel  <= 0;
    end else begin
        if( psg_cen     ) cnt<=cnt+1'd1;
        if( m2s_data    ) latch <= main_dout;
        if( psgdata_cs  ) psg_data <= dout;
        if( vlm_data_cs ) vlm_data <= dout;
        if( vlm_ctrl_cs ) { snd_en, vlm_rst, vlm_st, vlm_sel } <= A[8:3];
        if( rdac_cs     ) rdac <= dout;
    end
end

always @* begin
    rom_cs      = 0;
    ram_cs      = 0;
    latch_cs    = 0;
    cnt_cs      = 0;
    vlm_data_cs = 0;
    vlm_ctrl_cs = 0;
    rdac_cs     = 0;
    psgdata_cs  = 0;
    psg_cs      = 0;
    if( !mreq_n ) begin
        case(A[15:13])
            0,1: rom_cs    = 1;
            2: ram_cs      = 1; // 4000
            3: latch_cs    = 1; // 6000
            4: cnt_cs      = 1; // 8000
            5: vlm_data_cs = 1; // A000
            6: vlm_ctrl_cs = 1; // C000
            7: case( A[2:0] )
                0: rdac_cs    = 1;  // E000
                1: psgdata_cs = 1;  // E001
                2: psg_cs     = 1;  // E002
                default:;
            endcase
            default:;
        endcase
    end
end

always @(posedge clk) begin
    din  <= rom_cs   ? rom_data :
            ram_cs   ? ram_dout :
            cnt_cs   ? { 5'h1f, vlm_bsy, cnt[CNTW-1:CNTW-2] }  :
            latch_cs ? latch    :
            8'hff;
end

jt89 u_psg(
    .rst    ( rst           ),
    .clk    ( clk           ),
    .clk_en ( psg_cen       ),
    .wr_n   ( rdy1          ),
    .cs_n   ( ~psg_cs       ),
    .din    ( psg_data      ),
    .sound  ( psg_snd       ),
    .ready  ( rdy1          )
);

`ifndef VERILATOR
vlm5030_gl u_vlm(
    .i_rst   ( vlm_rst      ),
    .i_clk   ( clk          ),
    .i_oscen ( vlm_ceng     ),
    .i_start ( vlm_st       ),
    .i_vcu   ( 1'b0         ),
    .i_tst1  ( 1'b0         ),
    .o_tst2  (              ),
    .o_tst4  (              ),
    .i_d     ( vlm_mux      ),
    .o_a     ( { pcm_nc, pcm_addr[12:0] } ),
    .o_me_l  ( vlm_me_b     ),
    .o_mte   (              ),
    .o_bsy   ( vlm_bsy      ),

    .o_dao   (              ),
    .o_audio ( vlm_snd      )
);
`else
    reg busy_dummy=0;
    reg cnt_csl;

    assign vlm_bsy = busy_dummy;

    always @(posedge clk) begin
        cnt_csl <= cnt_cs;
        if( cnt_cs && !cnt_csl ) busy_dummy <= ~busy_dummy;
    end
`endif

wire signed [7:0] rdac_s;

jtframe_dcrm #(.SW(8)) u_dcrm(
    .rst    ( rst       ),
    .clk    ( clk       ),
    .sample ( cnt[6]    ),  // 14 kHz
    .din    ( rdac      ),
    .dout   ( rdac_s    )
);

wire [7:0] gain_psg  = !snd_en[2] ? 8'h18 : 8'h0;
wire [7:0] gain_vlm  = !snd_en[1] ? 8'h18 : 8'h0;
wire [7:0] gain_rdac = !snd_en[0] ? 8'h10 : 8'h0;

jtframe_mixer #(.W0(11),.W1(10),.W2(8)) u_mixer(
    .rst    ( rst       ),
    .clk    ( clk       ),
    .cen    ( psg_cen   ),
    // input signals
    .ch0    ( psg_snd   ),
    .ch1    ( vlm_snd   ),
    .ch2    ( rdac_s    ),
    .ch3    ( 16'd0     ),
    // gain for each channel in 4.4 fixed point format
    .gain0  ( gain_psg  ),
    .gain1  ( gain_vlm  ),
    .gain2  ( gain_rdac ),
    .gain3  ( 8'h00     ),
    .mixed  ( snd       ),
    .peak   ( peak      )
);

jtframe_ff u_irq(
    .rst      ( rst         ),
    .clk      ( clk         ),
    .cen      ( 1'b1        ),
    .din      ( 1'b1        ),
    .q        (             ),
    .qn       ( int_n       ),
    .set      (             ),
    .clr      ( irq_ack     ),
    .sigedge  ( m2s_on      )
);

/* verilator tracing_off */

jtframe_sysz80 #(.RAM_AW(10)) u_cpu(
    .rst_n      ( ~rst        ),
    .clk        ( clk         ),
    .cen        ( snd_cen     ),
    .cpu_cen    (             ),
    .int_n      ( int_n       ),
    .nmi_n      ( 1'b1        ),
    .busrq_n    ( 1'b1        ),
    .m1_n       ( m1_n        ),
    .mreq_n     ( mreq_n      ),
    .iorq_n     ( iorq_n      ),
    .rd_n       (             ),
    .wr_n       (             ),
    .rfsh_n     (             ),
    .halt_n     (             ),
    .busak_n    (             ),
    .A          ( A           ),
    .cpu_din    ( din         ),
    .cpu_dout   ( dout        ),
    .ram_dout   ( ram_dout    ),
    // manage access to ROM data from SDRAM
    .ram_cs     ( ram_cs      ),
    .rom_cs     ( rom_cs      ),
    .rom_ok     ( rom_ok      )
);

endmodule
